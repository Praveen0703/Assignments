`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.08.2025 14:23:50
// Design Name: 
// Module Name: question_13dt
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module question_13dt();
reg [3:0]
a= 4'b110x;

initial begin

if (a==4'b1100)
begin: B1 end
else
begin: B2 end
end
endmodule