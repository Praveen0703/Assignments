`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.08.2025 10:56:36
// Design Name: 
// Module Name: question_6dt
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test;
parameter WIDTH=8;

endmodule
module top;
test OUT ( ) ;
initial begin
OUT.WIDTH=10;
end
endmodule

