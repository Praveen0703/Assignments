`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.08.2025 12:37:44
// Design Name: 
// Module Name: question_12dt
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module question_12dt();
reg [3:0]a;
reg [6:0]b;
initial begin
a=4'd10;
b={a,1'b1};
end
endmodule
